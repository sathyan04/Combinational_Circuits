module encode_tb();
reg [3:0] in;
wire [1:0] out;
encode dut(.in(in),.out(out));
initial begin
	$monitor("Input=%b | Output=%b | Time=%0t",in,out,$time);
	$dumpfile("encodegtk.vcd");
	$dumpvars(0);
	in=4'b0000;#10;
	$display("");
	in=4'b0001;#10;
	$display("");
	in=4'b0010;#10;
	in=4'b0011;#10;
	$display("");
	in=4'b0100;#10;
	in=4'b0101;#10;
	in=4'b0110;#10;
	in=4'b0111;#10;
	$display("");
	in=4'b1000;#10;
	in=4'b1001;#10;
	in=4'b1010;#10;
	in=4'b1011;#10;
	in=4'b1100;#10;
	in=4'b1111;#10;
	in=4'b1110;#10;
	in=4'b1111;#10;
	$finish;
end
endmodule
